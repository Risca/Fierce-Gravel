../../src/FG_variables.vhd