../../src/FG_package.vhd